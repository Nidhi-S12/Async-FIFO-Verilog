module test;
  initial begin
    $display("FPGA Tools are working!");
    $finish;
  end
endmodule 